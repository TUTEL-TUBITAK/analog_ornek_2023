** sch_path: /home/ubuntu/Desktop/analog_ornek_2023/takim_adi_DTR/xschem/inv_TB.sch
**.subckt inv_TB
x1 A Y VDD GND inv
V1 VDD GND 1.8
V2 A GND pulse 0 1.8 2n 1n 1n 10n 20n
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt_mm





.control

save all

tran 0.1n 200n
save inv_TB.raw

.endc


**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/ubuntu/Desktop/analog_ornek_2023/takim_adi_DTR/xschem/inv.sym
** sch_path: /home/ubuntu/Desktop/analog_ornek_2023/takim_adi_DTR/xschem/inv.sch
.subckt inv  A Y VDD VSS
*.iopin A
*.iopin Y
*.iopin VDD
*.iopin VSS
XM1 Y A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
