* NGSPICE file created from inv_pex.ext - technology: sky130A

.subckt inv_pex A Y VDD VSS
X0 Y.t0 A.t0 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y.t1 A.t1 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
R0 A.n0 A.t1 485.228
R1 A.n0 A.t0 310.105
R2 A A.n0 0.963
R3 VSS.n6 VSS.n1 131.688
R4 VSS.n7 VSS.n6 93.294
R5 VSS.n18 VSS.t1 17.681
R6 VSS VSS.n18 0.303
R7 VSS.n16 VSS.n15 0.13
R8 VSS.n17 VSS.n16 0.13
R9 VSS.n18 VSS.n17 0.069
R10 VSS.n15 VSS.n8 0.015
R11 VSS.n8 VSS.n7 0.015
R12 VSS.n13 VSS.n12 0.007
R13 VSS.n12 VSS.n11 0.007
R14 VSS.n3 VSS.n2 0.003
R15 VSS.t0 VSS.n3 0.003
R16 VSS.n6 VSS.n5 0.003
R17 VSS.n13 VSS.n10 0.002
R18 VSS.n5 VSS.n4 0.002
R19 VSS.n10 VSS.n9 0.002
R20 VSS.n4 VSS.t0 0.001
R21 VSS.n1 VSS.n0 0.001
R22 VSS.n15 VSS.n14 0.001
R23 VSS.n14 VSS.n13 0.001
R24 Y.n0 Y.t0 18.864
R25 Y.n0 Y.t1 16.125
R26 Y Y.n0 0.177
R27 VDD.n12 VDD.n7 169.364
R28 VDD.n13 VDD.n12 105.135
R29 VDD.n18 VDD.t1 14.585
R30 VDD VDD.n18 0.486
R31 VDD.n16 VDD.n15 0.072
R32 VDD.n17 VDD.n16 0.072
R33 VDD.n18 VDD.n17 0.038
R34 VDD.n15 VDD.n14 0.006
R35 VDD.n14 VDD.n13 0.006
R36 VDD.n4 VDD.n1 0.003
R37 VDD.n1 VDD.n0 0.003
R38 VDD.n10 VDD.n9 0.003
R39 VDD.n12 VDD.n11 0.003
R40 VDD.n11 VDD.t0 0.003
R41 VDD.n9 VDD.n8 0.003
R42 VDD.n4 VDD.n3 0.001
R43 VDD.n3 VDD.n2 0.001
R44 VDD.t0 VDD.n10 0.001
R45 VDD.n15 VDD.n5 0.001
R46 VDD.n5 VDD.n4 0.001
R47 VDD.n7 VDD.n6 0.001
C0 VDD A 0.41fF
C1 VDD Y 1.25fF
C2 A Y 0.17fF
.ends

